library verilog;
use verilog.vl_types.all;
entity cod_vlg_vec_tst is
end cod_vlg_vec_tst;
