library verilog;
use verilog.vl_types.all;
entity vehi_vlg_vec_tst is
end vehi_vlg_vec_tst;
