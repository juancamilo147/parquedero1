library verilog;
use verilog.vl_types.all;
entity BCD7SEG_vlg_vec_tst is
end BCD7SEG_vlg_vec_tst;
