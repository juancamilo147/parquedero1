library verilog;
use verilog.vl_types.all;
entity cod is
    port(
        v               : in     vl_logic_vector(7 downto 0);
        f               : out    vl_logic_vector(3 downto 0)
    );
end cod;
